
VERSION             5.2 ;
NAMESCASESENSITIVE  ON ;
BUSBITCHARS         "()" ;
DIVIDERCHAR         "." ;


MACRO rf2_dec_bufad0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION INOUT ;
        PORT
            LAYER ALU2 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU2 ;
            RECT 24.00 29.00 26.00 31.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER ALU1 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
            RECT 4.00 9.00 6.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
    END
END rf2_dec_bufad0


MACRO rf2_dec_bufad1_l
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 19.00 31.00 21.00 ;
    END
END rf2_dec_bufad1_l


MACRO rf2_dec_bufad1_r
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END nq
    PIN q
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END q
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END i
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 98.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 19.00 31.00 21.00 ;
    END
END rf2_dec_bufad1_r


MACRO rf2_dec_bufad2_l
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      50.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq0
        DIRECTION INOUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END nq0
    PIN nq1
        DIRECTION INOUT ;
        PORT
            LAYER ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nq1
    PIN q0
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END q0
    PIN q1
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END q1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 47.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 47.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 48.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 19.00 46.00 21.00 ;
    END
END rf2_dec_bufad2_l


MACRO rf2_dec_bufad2_r
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      100.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq0
        DIRECTION INOUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END nq0
    PIN nq1
        DIRECTION INOUT ;
        PORT
            LAYER ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END nq1
    PIN q0
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 19.00 19.00 21.00 21.00 ;
        END
    END q0
    PIN q1
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END q1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 39.00 19.00 41.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 97.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 97.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 98.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 19.00 46.00 21.00 ;
    END
END rf2_dec_bufad2_r


MACRO rf2_dec_nand2
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i0
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 68.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 19.00 26.00 21.00 ;
        RECT 14.00 19.00 46.00 21.00 ;
    END
END rf2_dec_nand2


MACRO rf2_dec_nand3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 68.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 19.00 26.00 21.00 ;
        RECT 14.00 19.00 46.00 21.00 ;
    END
END rf2_dec_nand3


MACRO rf2_dec_nand4
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      70.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 44.00 19.00 46.00 21.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 19.00 26.00 21.00 ;
        END
    END i1
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 19.00 31.00 21.00 ;
        END
    END i2
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 14.00 19.00 16.00 21.00 ;
        END
    END i0
    PIN i3
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 34.00 19.00 36.00 21.00 ;
        END
    END i3
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 67.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 67.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 68.50 41.00 ;
        LAYER ALU2 ;
        RECT 14.00 19.00 46.00 21.00 ;
        RECT 19.00 19.00 26.00 21.00 ;
    END
END rf2_dec_nand4


MACRO rf2_dec_nao3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END nq
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i1
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 19.00 34.00 21.00 36.00 ;
        END
    END i2
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
        LAYER ALU2 ;
        RECT 4.00 19.00 11.00 21.00 ;
    END
END rf2_dec_nao3


MACRO rf2_dec_nbuf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      105.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
            RECT 14.00 9.00 16.00 11.00 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END nq
    PIN i
        DIRECTION INPUT ;
        PORT
            LAYER ALU1 ;
            RECT 49.00 39.00 51.00 41.00 ;
            RECT 49.00 34.00 51.00 36.00 ;
            RECT 49.00 29.00 51.00 31.00 ;
            RECT 49.00 24.00 51.00 26.00 ;
            RECT 49.00 19.00 51.00 21.00 ;
            RECT 49.00 14.00 51.00 16.00 ;
            RECT 49.00 9.00 51.00 11.00 ;
        END
    END i
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 102.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 102.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 103.50 41.00 ;
    END
END rf2_dec_nbuf


MACRO rf2_dec_nor3
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN nq
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU2 ;
            RECT 9.00 14.00 11.00 16.00 ;
        END
    END nq
    PIN i0
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 9.00 39.00 11.00 41.00 ;
        END
    END i0
    PIN i2
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END i2
    PIN i1
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 4.00 19.00 6.00 21.00 ;
        END
    END i1
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
        LAYER ALU2 ;
        RECT 4.00 19.00 11.00 21.00 ;
    END
END rf2_dec_nor3


MACRO rf2_inmux_buf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN sel0
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 34.00 39.00 36.00 41.00 ;
        END
    END sel0
    PIN sel1
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 14.00 26.00 16.00 ;
        END
    END sel1
    PIN sel
        DIRECTION INPUT ;
        PORT
            LAYER ALU1 ;
            RECT 14.00 89.00 16.00 91.00 ;
            RECT 14.00 84.00 16.00 86.00 ;
            RECT 14.00 79.00 16.00 81.00 ;
            RECT 14.00 74.00 16.00 76.00 ;
            RECT 14.00 69.00 16.00 71.00 ;
        END
    END sel
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 42.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 42.00 97.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
        RECT 1.50 59.00 43.50 91.00 ;
        LAYER ALU2 ;
        RECT 26.00 39.00 40.00 41.00 ;
        RECT 8.00 14.00 26.00 16.00 ;
        RECT 4.00 14.00 26.00 16.00 ;
        RECT 24.00 39.00 41.00 41.00 ;
    END
END rf2_inmux_buf


MACRO rf2_inmux_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      45.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN dinx
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU2 ;
            RECT 9.00 9.00 11.00 11.00 ;
        END
    END dinx
    PIN datain1
        DIRECTION INPUT ;
        PORT
            LAYER ALU1 ;
            RECT 39.00 39.00 41.00 41.00 ;
            RECT 39.00 34.00 41.00 36.00 ;
            RECT 39.00 29.00 41.00 31.00 ;
            RECT 39.00 24.00 41.00 26.00 ;
            RECT 39.00 19.00 41.00 21.00 ;
            RECT 39.00 14.00 41.00 16.00 ;
        END
    END datain1
    PIN datain0
        DIRECTION INPUT ;
        PORT
            LAYER ALU1 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END datain0
    PIN sel0
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 34.00 29.00 36.00 31.00 ;
        END
    END sel0
    PIN sel1
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 24.00 29.00 26.00 31.00 ;
        END
    END sel1
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 42.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 42.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 43.50 41.00 ;
        LAYER ALU2 ;
        RECT 24.00 29.00 36.00 31.00 ;
    END
END rf2_inmux_mem


MACRO rf2_mid_buf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN reada
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 19.00 59.00 21.00 61.00 ;
            RECT 19.00 54.00 21.00 56.00 ;
            RECT 19.00 49.00 21.00 51.00 ;
            RECT 19.00 44.00 21.00 46.00 ;
            RECT 19.00 39.00 21.00 41.00 ;
            RECT 19.00 34.00 21.00 36.00 ;
            RECT 19.00 29.00 21.00 31.00 ;
            RECT 19.00 24.00 21.00 26.00 ;
            RECT 19.00 19.00 21.00 21.00 ;
            RECT 19.00 14.00 21.00 16.00 ;
        END
    END reada
    PIN write
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 4.00 59.00 6.00 61.00 ;
            RECT 4.00 54.00 6.00 56.00 ;
            RECT 4.00 49.00 6.00 51.00 ;
            RECT 4.00 44.00 6.00 46.00 ;
            RECT 4.00 39.00 6.00 41.00 ;
            RECT 4.00 34.00 6.00 36.00 ;
            RECT 4.00 29.00 6.00 31.00 ;
            RECT 4.00 24.00 6.00 26.00 ;
            RECT 4.00 19.00 6.00 21.00 ;
            RECT 4.00 14.00 6.00 16.00 ;
        END
    END write
    PIN readb
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 59.00 31.00 61.00 ;
            RECT 29.00 54.00 31.00 56.00 ;
            RECT 29.00 49.00 31.00 51.00 ;
            RECT 29.00 44.00 31.00 46.00 ;
            RECT 29.00 39.00 31.00 41.00 ;
            RECT 29.00 34.00 31.00 36.00 ;
            RECT 29.00 29.00 31.00 31.00 ;
            RECT 29.00 24.00 31.00 26.00 ;
            RECT 29.00 19.00 31.00 21.00 ;
            RECT 29.00 14.00 31.00 16.00 ;
        END
    END readb
    PIN selrb
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 24.00 84.00 26.00 86.00 ;
        END
    END selrb
    PIN selra
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 14.00 84.00 16.00 86.00 ;
        END
    END selra
    PIN nck
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT -1.00 89.00 1.00 91.00 ;
        END
    END nck
    PIN selw
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 9.00 84.00 11.00 86.00 ;
        END
    END selw
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 32.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 32.00 97.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
        RECT 1.50 59.00 33.50 91.00 ;
        LAYER ALU2 ;
        RECT 14.00 64.00 31.00 66.00 ;
        RECT 4.00 59.00 31.00 61.00 ;
        RECT 4.00 39.00 31.00 41.00 ;
        RECT 14.00 19.00 26.00 21.00 ;
        RECT 4.00 14.00 31.00 16.00 ;
        RECT 17.00 39.00 21.00 41.00 ;
        RECT 17.00 14.00 21.00 16.00 ;
        RECT 14.00 64.00 21.00 66.00 ;
        RECT 24.00 64.00 31.00 66.00 ;
        LAYER ALU3 ;
        RECT 14.00 19.00 16.00 66.00 ;
        RECT 24.00 19.00 26.00 66.00 ;
        RECT 24.00 19.00 26.00 66.00 ;
        RECT 14.00 19.00 16.00 66.00 ;
    END
END rf2_mid_buf


MACRO rf2_mid_mem_r0
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN busb
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER ALU2 ;
            RECT 34.00 24.00 36.00 26.00 ;
        END
    END busb
    PIN busa
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER ALU2 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END busa
    PIN write
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END write
    PIN dinx
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END dinx
    PIN reada
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END reada
    PIN readb
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 29.00 31.00 31.00 ;
        END
    END readb
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 29.00 26.00 31.00 ;
    END
END rf2_mid_mem_r0


MACRO rf2_mid_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      35.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN busb
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER ALU2 ;
            RECT 34.00 24.00 36.00 26.00 ;
        END
    END busb
    PIN busa
        DIRECTION OUTPUT TRISTATE ;
        PORT
            LAYER ALU2 ;
            RECT 34.00 14.00 36.00 16.00 ;
        END
    END busa
    PIN write
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 4.00 29.00 6.00 31.00 ;
        END
    END write
    PIN dinx
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 19.00 9.00 21.00 11.00 ;
        END
    END dinx
    PIN reada
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 19.00 29.00 21.00 31.00 ;
        END
    END reada
    PIN readb
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 29.00 29.00 31.00 31.00 ;
        END
    END readb
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 32.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 32.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 33.50 41.00 ;
        LAYER ALU2 ;
        RECT 19.00 29.00 26.00 31.00 ;
        RECT 4.00 29.00 16.00 31.00 ;
    END
END rf2_mid_mem


MACRO rf2_out_buf
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      105.00 BY 100.00 ;
    SYMMETRY  Y ;
    SITE      core ;
    PIN xcks
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU3 ;
            RECT 14.00 59.00 16.00 61.00 ;
            RECT 14.00 54.00 16.00 56.00 ;
            RECT 14.00 49.00 16.00 51.00 ;
            RECT 14.00 44.00 16.00 46.00 ;
            RECT 14.00 39.00 16.00 41.00 ;
            RECT 14.00 34.00 16.00 36.00 ;
            RECT 14.00 29.00 16.00 31.00 ;
            RECT 14.00 24.00 16.00 26.00 ;
            RECT 14.00 19.00 16.00 21.00 ;
            RECT 14.00 14.00 16.00 16.00 ;
        END
    END xcks
    PIN nck
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU2 ;
            RECT 79.00 89.00 81.00 91.00 ;
            RECT 74.00 89.00 76.00 91.00 ;
            RECT 69.00 89.00 71.00 91.00 ;
            RECT 64.00 89.00 66.00 91.00 ;
            RECT 59.00 89.00 61.00 91.00 ;
            RECT 54.00 89.00 56.00 91.00 ;
            RECT 49.00 89.00 51.00 91.00 ;
            RECT 44.00 89.00 46.00 91.00 ;
            RECT 39.00 89.00 41.00 91.00 ;
            RECT 34.00 89.00 36.00 91.00 ;
            RECT 29.00 89.00 31.00 91.00 ;
            RECT 24.00 89.00 26.00 91.00 ;
            RECT 19.00 89.00 21.00 91.00 ;
            RECT 14.00 89.00 16.00 91.00 ;
            LAYER ALU2 ;
            RECT 14.00 89.00 16.00 91.00 ;
        END
    END nck
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 102.00 47.00 ;
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 53.00 102.00 53.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 102.00 3.00 ;
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 97.00 102.00 97.00 ;
        END
    END vss
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
            LAYER ALU1 ;
            RECT 99.00 89.00 101.00 91.00 ;
            RECT 99.00 84.00 101.00 86.00 ;
            RECT 99.00 79.00 101.00 81.00 ;
            RECT 99.00 74.00 101.00 76.00 ;
            RECT 99.00 69.00 101.00 71.00 ;
            RECT 99.00 64.00 101.00 66.00 ;
            RECT 99.00 59.00 101.00 61.00 ;
        END
    END ck
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 103.50 41.00 ;
        RECT 1.50 59.00 103.50 91.00 ;
        LAYER ALU2 ;
        RECT 9.00 59.00 21.00 61.00 ;
        RECT 9.00 39.00 21.00 41.00 ;
        RECT 9.00 14.00 21.00 16.00 ;
    END
END rf2_out_buf


MACRO rf2_out_mem
    CLASS     CORE ;
    ORIGIN    0.00 0.00 ;
    SIZE      105.00 BY 50.00 ;
    SYMMETRY  X Y ;
    SITE      core ;
    PIN dataoutb
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU1 ;
            RECT 44.00 39.00 46.00 41.00 ;
            RECT 44.00 34.00 46.00 36.00 ;
            RECT 44.00 29.00 46.00 31.00 ;
            RECT 44.00 24.00 46.00 26.00 ;
            RECT 44.00 19.00 46.00 21.00 ;
            RECT 44.00 14.00 46.00 16.00 ;
            RECT 44.00 9.00 46.00 11.00 ;
        END
    END dataoutb
    PIN dataouta
        DIRECTION OUTPUT ;
        PORT
            LAYER ALU1 ;
            RECT 59.00 39.00 61.00 41.00 ;
            RECT 59.00 34.00 61.00 36.00 ;
            RECT 59.00 29.00 61.00 31.00 ;
            RECT 59.00 24.00 61.00 26.00 ;
            RECT 59.00 19.00 61.00 21.00 ;
            RECT 59.00 14.00 61.00 16.00 ;
            RECT 59.00 9.00 61.00 11.00 ;
        END
    END dataouta
    PIN busb
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 4.00 24.00 6.00 26.00 ;
        END
    END busb
    PIN xcks
        DIRECTION INPUT ;
        PORT
            LAYER ALU3 ;
            RECT 14.00 24.00 16.00 26.00 ;
        END
    END xcks
    PIN busa
        DIRECTION INPUT ;
        PORT
            LAYER ALU2 ;
            RECT 99.00 14.00 101.00 16.00 ;
        END
    END busa
    PIN vdd
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 47.00 102.00 47.00 ;
        END
    END vdd
    PIN vss
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
            LAYER ALU1 ;
            WIDTH 6.00 ;
            PATH 3.00 3.00 102.00 3.00 ;
        END
    END vss
    OBS
        LAYER ALU1 ;
        RECT 1.50 9.00 103.50 41.00 ;
        LAYER ALU2 ;
        RECT 14.00 24.00 86.00 26.00 ;
        RECT 14.00 24.00 86.00 26.00 ;
    END
END rf2_out_mem


END LIBRARY
